library verilog;
use verilog.vl_types.all;
entity CPU289_vlg_vec_tst is
end CPU289_vlg_vec_tst;
