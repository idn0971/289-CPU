library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CPU289 is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity CPU289;

architecture RTL of CPU289 is

begin

end architecture RTL;
